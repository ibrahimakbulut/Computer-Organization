module mips32_single_cycle(clk,last_result);

wire [31:0] instruction;
input clk;
output [31:0] last_result;
wire [31:0] result;

wire [2:0] selects_bits_alue;
wire [31:0] rs,rt;
wire [31:0] dataA,dataB,shamt,result_sltu,result_temp;
wire [31:0] PC;
wire [31:0] immediate_extended_sign,immediate_extended_zero,result_immediate_extended;
wire [4:0] write_register;

wire reg_des,branch_signal,jump_signal,memread,memwrite,memtoreg,regwrite,alusrc;
wire temp_branch_signal;
wire or1,or2,or3,or4,or5;
wire[31:0] memory_data;
wire outbit,sltu_signal,zero_or_sign;

wire r_type_not,r_type;

wire[31:0] bus_b,bus_a,bus_b2;

wire [31:0] sub_equal;

or o11(r_type_not,instruction[31],instruction[30],instruction[29],instruction[28],instruction[27],instruction[26]);

not n8(r_type,r_type_not);  //instruction r type or not



full_minus_32 y5(rs,rt,1'b0,sub_equal,outbit);
or o1(or1,sub_equal[0],sub_equal[1],sub_equal[2],sub_equal[3],sub_equal[4],sub_equal[5],sub_equal[6],sub_equal[7],sub_equal[8]);
or o2(or2,sub_equal[9],sub_equal[10],sub_equal[11],sub_equal[12],sub_equal[13],sub_equal[14],sub_equal[15],sub_equal[16]);
or o3(or3,sub_equal[17],sub_equal[18],sub_equal[19],sub_equal[20],sub_equal[21],sub_equal[22],sub_equal[23],sub_equal[24]);
or o4(or4,sub_equal[25],sub_equal[26],sub_equal[27],sub_equal[28],sub_equal[29],sub_equal[30],sub_equal[31]);
or o5(or5,or4,or3,or2,or1);


//to call right operation control_unit function is called then selects bits are generated by it.
control_unit c1(selects_bits_alue,instruction[5:0],instruction[31:26],reg_des,branch_signal,jump_signal,memread,memwrite,memtoreg,regwrite,alusrc,zero_or_sign);

not n1(equal,or5);

and a1(temp_branch_signal,equal,branch_signal);

next_PC v1(temp_branch_signal,jump_signal,clk,instruction[31:0],PC);

instruction_memory v2(PC,instruction,clk);

//rt or rd is chosen as a write register
mux5_2_1 m0(reg_des,instruction[20:16],instruction[15:11],write_register);

//call the mips_register function
mips_registers f1(rs,rt,last_result,instruction[25:21],instruction[20:16],write_register,1'b1,clk);


buf h1(shamt[0],instruction[6]);
buf h2(shamt[1],instruction[7]);
buf h3(shamt[2],instruction[8]);
buf h4(shamt[3],instruction[9]);
buf h5(shamt[4],instruction[10]);
buf h6(shamt[5],1'b0);
buf h7(shamt[6],1'b0);
buf h8(shamt[7],1'b0);
buf h9(shamt[8],1'b0); //shift amount is assigned to shamt wire.
buf h10(shamt[9],1'b0);
buf h11(shamt[10],1'b0);
buf h12(shamt[11],1'b0);
buf h13(shamt[12],1'b0);
buf h14(shamt[13],1'b0);
buf h15(shamt[14],1'b0);
buf h16(shamt[15],1'b0);
buf h17(shamt[16],1'b0);
buf h18(shamt[17],1'b0);
buf h19(shamt[18],1'b0);
buf h20(shamt[19],1'b0);
buf h21(shamt[20],1'b0);
buf h22(shamt[21],1'b0);
buf h23(shamt[22],1'b0);
buf h24(shamt[23],1'b0);
buf h25(shamt[24],1'b0);
buf h26(shamt[25],1'b0);
buf h27(shamt[26],1'b0);
buf h28(shamt[27],1'b0);
buf h29(shamt[28],1'b0);
buf h30(shamt[29],1'b0);
buf h31(shamt[30],1'b0);
buf h32(shamt[31],1'b0);

sign_extender p1(instruction[15:0],immediate_extended_sign);
zero_extender p2(instruction[15:0],immediate_extended_zero);

//immediate zero extended or sign extended choisen
mux32_2_1 m45(zero_or_sign,immediate_extended_sign,immediate_extended_zero,result_immediate_extended);

//if operation shift then rt must be choisen instead of rs,shamt must be choisen instead of rt.
mux32_2_1 m1(instruction[5],rt,rs,dataA);
mux32_2_1 m2(instruction[5],shamt,rt,dataB);

mux32_2_1 m3(alusrc,dataB,result_immediate_extended,bus_b);
mux32_2_1 m8(r_type,rs,dataA,bus_a);

//operation is performed after selecting the datas
alu32 a2(bus_a,bus_b,selects_bits_alue,result_temp);

mux32_2_1 m9(r_type,rt,dataB,bus_b2);
data_memory t1(result,bus_b2,memory_data,memwrite,memread,clk);

mux32_2_1 m5(memtoreg,result,memory_data,last_result);

//The most important bit of the alu32 result is combined with the result_sltu
buf d1(result_sltu[0],result_temp[31]);
buf d2(result_sltu[1],1'b0);
buf d3(result_sltu[2],1'b0);
buf d4(result_sltu[3],1'b0);
buf d5(result_sltu[4],1'b0);
buf d6(result_sltu[5],1'b0);
buf d7(result_sltu[6],1'b0);
buf d8(result_sltu[7],1'b0);
buf d9(result_sltu[8],1'b0);
buf d10(result_sltu[9],1'b0);
buf d11(result_sltu[10],1'b0);  
buf d12(result_sltu[11],1'b0);
buf d13(result_sltu[12],1'b0);
buf d14(result_sltu[13],1'b0);
buf d15(result_sltu[14],1'b0);
buf d16(result_sltu[15],1'b0);
buf d17(result_sltu[16],1'b0);
buf d18(result_sltu[17],1'b0);
buf d19(result_sltu[18],1'b0);
buf d20(result_sltu[19],1'b0);
buf d21(result_sltu[20],1'b0);
buf d22(result_sltu[21],1'b0);
buf d23(result_sltu[22],1'b0);
buf d24(result_sltu[23],1'b0);
buf d25(result_sltu[24],1'b0);
buf d26(result_sltu[25],1'b0);
buf d27(result_sltu[26],1'b0);
buf d28(result_sltu[27],1'b0);
buf d29(result_sltu[28],1'b0);
buf d30(result_sltu[29],1'b0);
buf d31(result_sltu[30],1'b0);
buf d32(result_sltu[31],1'b0);

and a45(sltu_signal,r_type,instruction[3]);

//If the operation is sltu then chosen the result_sltu ,if not chosen result_temp(which is result of alu32)
mux32_2_1 m4(sltu_signal,result_temp,result_sltu,result);

endmodule