
module alu32_testbench(); 
reg [31:0] in1, in2;
wire [31:0] result;
reg [2:0] select;


alu32 alu_test(in1,in2,select,result);

initial begin
in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; select = 3'b000;  
#50;
in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; select = 3'b001;  
#50;
in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; select = 3'b010;  
#50;
in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; select = 3'b011;  
#50;
in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; select = 3'b100;  
#50;
in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; select = 3'b101;  
#50;
in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; select = 3'b110;  
#50;
in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; select = 3'b111; 
#50;



in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; select = 3'b000;
#50;
in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; select = 3'b001;
#50;
in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; select = 3'b010;
#50;
in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; select = 3'b011;
#50;
in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; select = 3'b100;
#50;
in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; select = 3'b101;
#50;
in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; select = 3'b110;
#50;
in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; select = 3'b111;
#50;


in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; select = 3'b000;
#50;
in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; select = 3'b001;
#50;
in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; select = 3'b010;
#50;
in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; select = 3'b011;
#50;
in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; select = 3'b100;
#50;
in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; select = 3'b101;
#50;
in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; select = 3'b110;
#50;
in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; select = 3'b111;
#50;
end
 
 
initial
begin
$monitor("time = %2d, in1 = %32b, in2= %32b, opcode= %3b, result = %32b \n" , $time, in1, in2,select,result);
end
 
 
 endmodule